//PWM Controller SystemVerilog description

module pwm
  #(PARAMETER FREQ = 100)
   (input logic [7:0] duty_cycle,
    output logic out);

   pipo_reg dc(


endmodule: pwm
